LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MEMORIA IS
	PORT(CLK, RST, WR : IN STD_LOGIC;
			ADDRESS: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_IN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_IN_00, P_IN_01, P_IN_02, P_IN_03 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_IN_04, P_IN_05, P_IN_06, P_IN_07 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_IN_08, P_IN_09, P_IN_10, P_IN_11 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_IN_12, P_IN_13, P_IN_14, P_IN_15 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_00, P_OUT_01, P_OUT_02, P_OUT_03 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_04, P_OUT_05, P_OUT_06, P_OUT_07 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_08, P_OUT_09, P_OUT_10, P_OUT_11 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_12, P_OUT_13, P_OUT_14, P_OUT_15 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END ENTITY;
	
	
	ARCHITECTURE RTL OF MEMORIA IS
		COMPONENT mem_programa IS
			PORT(CLK: IN STD_LOGIC;
			ADDREES: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
			
		END COMPONENT mem_programa;
		
		
		COMPONENT mem_datos IS
			PORT(CLK, WR: IN STD_LOGIC;
			ADDREES: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			DATA_IN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
			
		END COMPONENT mem_datos;
		
		
		COMPONENT puertos_salida IS

			PORT(	CLK, RST, WR: IN STD_LOGIC;
			ADDRESS     : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA_IN     : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_00, P_OUT_01, P_OUT_02, P_OUT_03: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_04, P_OUT_05, P_OUT_06, P_OUT_07: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_08, P_OUT_09, P_OUT_10, P_OUT_11: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			P_OUT_12, P_OUT_13, P_OUT_14, P_OUT_15: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
		END COMPONENT puertos_salida;
		
		SIGNAL ROM_OUT, RAM_OUT: STD_LOGIC_VECTOR(7 downto 0);
		SIGNAL OUTPUT_PORT_ADDR: STD_LOGIC_VECTOR(3 DOWNTO 0);
		SIGNAL RAM_ADDRESS, ROM_ADDRESS: STD_LOGIC_VECTOR(6 DOWNTO 0);
		
		
		BEGIN
			ROM_ADDRESS <= ADDRESS(6 DOWNTO 0) WHEN (ADDRESS(7) = '0') ELSE "0000000";
			RAM_ADDRESS <= ADDRESS(6 DOWNTO 0) WHEN (ADDRESS(7) = '0') ELSE "0000000";
			OUTPUT_PORT_ADDR <= ADDRESS(3 DOWNTO 0) WHEN (ADDRESS(7 DOWNTO 4)= X"F") ELSE "0000";
			
			MEM_PROG : mem_programa port map(CLK, ROM_ADDRESS, ROM_OUT);
			MEM_DAT  : mem_datos port map(CLK, WR, RAM_ADDRESS, DATA_IN, RAM_OUT);
			PUERTOS  : PUErtos_salida port map(CLK, RST, WR, OUTPUT_PORT_ADDR, DATA_IN, P_OUT_00,P_OUT_01,P_OUT_02, P_OUT_03,
																	P_OUT_04, P_OUT_05, P_OUT_06, P_OUT_07, P_OUT_08, P_OUT_09, P_OUT_10, P_OUT_11,
																	P_OUT_12, P_OUT_13, P_OUT_14, P_OUT_15);
																	
			
			DATA_OUT <= ROM_OUT WHEN ADDRESS < X"80" ELSE
							RAM_OUT WHEN ADDRESS < X"E0" ELSE
							P_IN_00 WHEN ADDRESS = X"F0" ELSE
							P_IN_01 WHEN ADDRESS = X"F1" ELSE
							P_IN_02 WHEN ADDRESS = X"F2" ELSE
							P_IN_03 WHEN ADDRESS = X"F3" ELSE
							P_IN_04 WHEN ADDRESS = X"F4" ELSE
							P_IN_05 WHEN ADDRESS = X"F5" ELSE
							P_IN_06 WHEN ADDRESS = X"F6" ELSE
							P_IN_07 WHEN ADDRESS = X"F7" ELSE
							P_IN_08 WHEN ADDRESS = X"F8" ELSE
							P_IN_09 WHEN ADDRESS = X"F9" ELSE
							P_IN_10 WHEN ADDRESS = X"FA" ELSE
							P_IN_11 WHEN ADDRESS = X"FB" ELSE
							P_IN_12 WHEN ADDRESS = X"FC" ELSE
							P_IN_13 WHEN ADDRESS = X"FD" ELSE
							P_IN_14 WHEN ADDRESS = X"FE" ELSE
							P_IN_15 WHEN ADDRESS = X"FF" ELSE
							X"00";
			END ARCHITECTURE;
							
							

			
		
		
		
		
		
		
		
		
		
		
		
		
		