LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY mem_programa IS
	 PORT(CLK: IN STD_LOGIC;
			ADDREES: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			DATA_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
			
	END mem_programa;
	
	
ARCHITECTURE RTL OF mem_programa IS

	CONSTANT LDA_INM: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"86";
	CONSTANT LDB_INM: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"87";
	CONSTANT LDA_DIR: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"88";
	CONSTANT LDB_DIR: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"89";
	CONSTANT STORE_A: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"96";
	CONSTANT STORE_B: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"97";

	
	
	CONSTANT ADD_AB: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"40";
	CONSTANT SUB_AB: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"41";
	CONSTANT AND_AB: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"42";
	CONSTANT OR_AB: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"43";
	CONSTANT XOR_AB: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"44";
	CONSTANT INC_A: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"45";
	CONSTANT INC_B: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"46";
	CONSTANT DEC_A: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"47";
	CONSTANT DEC_B: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"48";
	CONSTANT NOT_A: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"50";
	CONSTANT NOT_B: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"51";
	
	
	
	CONSTANT JMP: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"20";
	CONSTANT JN: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"21";
	CONSTANT JNN: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"22";
	CONSTANT JZ: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"23";
	CONSTANT JNZ: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"24";
	CONSTANT JOV: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"25";
	CONSTANT JNOV: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"26";
	CONSTANT JC: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"27";
	CONSTANT JNC: STD_LOGIC_VECTOR(7 DOWNTO 0) := X"28";
	
	TYPE instmem is ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	SIGNAL ROM: instmem :=( 0    =>  LDA_DIR,
									1    =>  X"F0",
									2    => LDB_DIR,
									3    => X"F1",
									4    => STORE_A,
									5    => X"E3",
									6    => STORE_B,
									7    => X"E3",
									8    => ADD_AB,
									9    => STORE_A,
									10    => X"E3",
									
									
									
									
									
									
									OTHERS => X"00");
									
									
	BEGIN
		PROCESS(CLK)
			BEGIN
				IF(CLK' EVENT AND CLK = '1') THEN
					DATA_OUT <= ROM(CONV_INTEGER(UNSIGNED(ADDREES)));
				END IF;
			END PROCESS;
	END ARCHITECTURE;
	

			