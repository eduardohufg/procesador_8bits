LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY BIT_SLICE IS

	PORT ( A,B: IN STD_LOGIC;
			NA,NB,CIN: IN STD_LOGIC;
			AANDB, NEGB, NEGA, AXORB, AORB, AMASB: IN STD_LOGIC;
			C, S: OUT STD_LOGIC
	);
	
END BIT_SLICE;

ARCHITECTURE RTL OF BIT_SLICE IS

	COMPONENT ha IS

		PORT (a,b : IN STD_LOGIC;
      s, Cout: OUT STD_LOGIC);
	END COMPONENT ha;
	
	SIGNAL XORAIN, XORBIN: STD_LOGIC;
	SIGNAL ORINTCONT: STD_LOGIC;
	SIGNAL COUTHA1: STD_LOGIC;
	SIGNAL SOUTHA1: STD_LOGIC;
	SIGNAL COUTHA2: STD_LOGIC;
	SIGNAL SOUTHA2: STD_LOGIC;

	SIGNAL AND1: STD_LOGIC;
	SIGNAL AND2: STD_LOGIC;
	SIGNAL AND3: STD_LOGIC;
	SIGNAL AND4: STD_LOGIC;
	SIGNAL AND5: STD_LOGIC;
	SIGNAL OR1: STD_LOGIC;
	SIGNAL ANDAUX: STD_LOGIC;
	SIGNAL ORGRAND: STD_LOGIC;
	SIGNAL SOUT: STD_LOGIC;
	
	BEGIN
	
	XORAIN <= A XOR NA;
	XORBIN <= B XOR NB;
	ORINTCONT <= NA OR NB OR CIN;
	
	I0: ha PORT MAP(XORAIN, XORBIN, SOUTHA1, COUTHA1);
	I1: ha PORT MAP(SOUTHA1, ORINTCONT, SOUTHA2, COUTHA2);
	
	C <= COUTHA1 OR COUTHA2;
	
	AND1 <= COUTHA1 AND AANDB;
	AND2 <= XORBIN AND NEGB;
	AND3 <= XORAIN AND NEGA;
	AND4 <= SOUTHA1 AND AXORB;
	AND5 <= SOUTHA2 AND AMASB;
	OR1 <= XORAIN OR XORBIN;
	ANDAUX <= OR1 AND AORB;
	ORGRAND <= AND1 OR AND2 OR AND3 OR ANDAUX OR AND4;
	S <= ORGRAND OR AND5;
	
	
	
	END RTL;
	
	
	